LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
ENTITY REG_Test IS
END REG_Test;
 
ARCHITECTURE behavior OF REG_Test IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT REG
    PORT(
         I_REG_EN : IN  std_logic;
         I_REG_WE : IN  std_logic;
         I_REG_SEL_RS : IN  std_logic_vector(4 downto 0);
         I_REG_SEL_RT : IN  std_logic_vector(4 downto 0);
         I_REG_SEL_RD : IN  std_logic_vector(4 downto 0);
         I_REG_DATA_RD : IN  std_logic_vector(31 downto 0);
         O_REG_DATA_A : OUT  std_logic_vector(31 downto 0);
         O_REG_DATA_B : OUT  std_logic_vector(31 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal I_REG_EN : std_logic := '0';
   signal I_REG_WE : std_logic := '0';
   signal I_REG_SEL_RS : std_logic_vector(4 downto 0) := (others => '0');
   signal I_REG_SEL_RT : std_logic_vector(4 downto 0) := (others => '0');
   signal I_REG_SEL_RD : std_logic_vector(4 downto 0) := (others => '0');
   signal I_REG_DATA_RD : std_logic_vector(31 downto 0) := (others => '0');

 	--Outputs
   signal O_REG_DATA_A : std_logic_vector(31 downto 0);
   signal O_REG_DATA_B : std_logic_vector(31 downto 0);
   -- No clocks detected in port list. Replace <clock> below with 
   -- appropriate port name 
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: REG PORT MAP (
          I_REG_EN => I_REG_EN,
          I_REG_WE => I_REG_WE,
          I_REG_SEL_RS => I_REG_SEL_RS,
          I_REG_SEL_RT => I_REG_SEL_RT,
          I_REG_SEL_RD => I_REG_SEL_RD,
          I_REG_DATA_RD => I_REG_DATA_RD,
          O_REG_DATA_A => O_REG_DATA_A,
          O_REG_DATA_B => O_REG_DATA_B
        );

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	

      -- insert stimulus here 
		I_REG_EN <= '1';
		I_REG_SEL_RS <= "00000";
		I_REG_SEL_RT <= "00010";
		wait for 20 ns;
		
		I_REG_SEL_RS <= "01010";
		I_REG_SEL_RT <= "01011";
		wait for 20 ns;
		
		I_REG_WE <= '1';
		I_REG_SEL_RD <= "01010";
		I_REG_DATA_RD <= x"FFFFFFFF";
		wait for 20 ns;
		
		I_REG_WE <= '0';
      wait for 20 ns;
		
		I_REG_WE <= '1';
		I_REG_SEL_RD <= "01011";
		I_REG_DATA_RD <= x"AAAAAAAA";
		wait for 20 ns;
		
		I_REG_WE <= '0';
      wait;
   end process;

END;
